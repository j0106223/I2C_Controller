module i2c_mem_model (

);
    input clk;
    input reset_n;
    
    input scl;
    input sda;
    output scl;
    output sda;

endmodule 