module i2c_core (
    
);
endmodule